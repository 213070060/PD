`timescale 1ns / 1ps
module testbench;  
	reg clk;  
	reg reset;   
	wire [15:0] pc_out;  
	wire [15:0] alu_result;
	integer i;
	processor uut (.clk(clk), .reset(reset), .pc_out(pc_out), .alu_result(alu_result));  
	initial begin  
		clk = 0;  
		for (i=0;i<=100;i = i+1) begin
			#10 clk = ~clk;
		end
	end  
	initial begin 
		reset = 1;
		#100; // Wait 100 ns for global reset to finish
		reset = 0; 
		// Add stimulus here  
	end  
endmodule