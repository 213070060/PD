module instr_mem (  
      input     [15:0]     pc,  
      output wire     [15:0]          instruction );  
      
	  wire [4 : 0] rom_addr = pc[5 : 1];  
      reg [15:0] rom[31:0];  
								 //Sa  Sb  Dest
      initial begin  			 //Ra  Rb  Rc	
				rom[0]  = 16'b0001_001_010_011_0_00; // add R3 = R1 + R2 = 5
				rom[1]  = 16'b0001_000_011_101_0_10; // adc R5 = R3 + R0 = no change since cy = 0
				rom[2]  = 16'b0000_110_100_111111; //adi R4 = R6+FFFF = 6, cy = 1 
				rom[3]  = 16'b0001_010_011_101_0_10; //adc R5 = R3+R2 = 8
				rom[4]  = 16'b0001_000_011_101_0_01; //adz R5 = R0 + R3 = no change if z=1 (R5 - no change) 
				rom[5]  = 16'b0000_000_101_111111; //adi R5 = R0 +FFFF = 0, z = 1 
				rom[6]  = 16'b0001_000_011_101_0_01; //adz R5 = R0+R3 = 6 
				rom[7]  = 16'b0010_000_010_110_0_00; //ndu R6= R0 nand R2 = FFFE 
				rom[8]  = 16'b0000_000_101_111111; //adi R5 = R0 + FFFF = 0, z =1
				rom[9]  = 16'b0010_000_011_101_0_01; //ndz R5 = R0 nand R3 = FFFE
				rom[10] = 16'b0000_000_110_111111; // adi R6 = R0 + FFFF = 0, c = z =1 
				rom[11] = 16'b0010_010_011_101_0_10; //ndc  R5 = R3 nand R2 = FFFE 
				rom[12] = 16'b0001_000_001_101_0_11; //adl R5 = <<R1 + R0 = 5 
				rom[13] = 16'b0000_001_000_000001; //adi R0 = R1 + 1 = 3
				rom[14] = 16'b0011_101_000_000_111; // lhi R5 = 0380
				rom[15] = 16'b0101_010_110_000001; //sw mem(R6+1) = R2 = 3
				rom[16] = 16'b0100_101_110_000_001; //lw R5 = mem(8) = 3
				rom[17] = 16'b1000_000_010_000101; //BEQ PC<=change to 2e
				rom[18] = 16'b0000_000_000_000000; //nop
				rom[19] = 16'b0000_000_000_000000; //nop
				rom[20] = 16'b0000_000_000_000000; //nop
				rom[21] = 16'b0000_000_000_000000; //nop
				rom[22] = 16'b0000_000_000_000000; //nop
				rom[23] = 16'b1001_101_000000100; //JAL PC<=PC+0100<=27
				rom[24] = 16'b1000_000_010_000010; //BEQ PC<=PC+2<=22 since R0=R2=3
				rom[19] = 16'b0000_000_000_000000; //nop
				rom[20] = 16'b0000_000_000_000000; //nop
				rom[21] = 16'b0000_000_000_000000; //nop
				rom[22] = 16'b0000_000_101_011010; //adi R5 = R4+20 = 26
				rom[23] = 16'b1010_000_101_000000; //JLR R0 R5
				rom[24] = 16'b0000_000_000_000000; //nop
				rom[25] = 16'b0000_000_000_000000; //nop
				rom[26] = 16'b1011_000_000_011010; //JRI PC<=R2+26 = 38
				rom[27] = 16'b0000_000_000_000000; //nop
				rom[28] = 16'b0000_000_000_000000; //nop
				rom[29] = 16'b0000_000_000_000000; //nop
				rom[30] = 16'b0000_000_000_000000; //nop
				rom[31] = 16'b0000_000_000_000000; //nop

     end  
     assign instruction = (pc[15:0] < 64 )? rom[rom_addr[4:0]]: 16'd0;  
 endmodule   
